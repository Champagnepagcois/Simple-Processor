module bit_register ( 
	clk,
	reset,
	data_in,
	data_out
	) ;

input  clk;
input  reset;
input  data_in;
inout  data_out;
